module Forward(

	//MODULE INPUTS



	//MODULE OUTPUTS



);

endmodule
