module Forward(

	//MODULE INPUTS
		input [4:0] ID/EX.RegisterRt,
		input [4:0] ID/EX.RegisterRs,
		input [4:0] MEM/WB.RegisterRd,
		input EX/MEM.RegWrite,
		input MEM/WB.RegWrite,

	//MODULE OUTPUTS
		output [1:0] ForwardA,
		output [1:0] ForwardB



);

endmodule
